
module CU(clk, bus);
	input wire clk;
	inout wire[15:0] bus;

endmodule

module register ( index, bus, rEn, wEn, reset );
  input [3:0] index;
  inout [15:0] bus;
  input rEn, wEn, reset;
  wire   \register[3][15] , \register[3][14] , \register[3][13] ,
         \register[3][12] , \register[3][11] , \register[3][10] ,
         \register[3][9] , \register[3][8] , \register[3][7] ,
         \register[3][6] , \register[3][5] , \register[3][4] ,
         \register[3][3] , \register[3][2] , \register[3][1] ,
         \register[3][0] , \register[2][15] , \register[2][14] ,
         \register[2][13] , \register[2][12] , \register[2][11] ,
         \register[2][10] , \register[2][9] , \register[2][8] ,
         \register[2][7] , \register[2][6] , \register[2][5] ,
         \register[2][4] , \register[2][3] , \register[2][2] ,
         \register[2][1] , \register[2][0] , \register[1][15] ,
         \register[1][14] , \register[1][13] , \register[1][12] ,
         \register[1][11] , \register[1][10] , \register[1][9] ,
         \register[1][8] , \register[1][7] , \register[1][6] ,
         \register[1][5] , \register[1][4] , \register[1][3] ,
         \register[1][2] , \register[1][1] , \register[1][0] ,
         \register[0][15] , \register[0][14] , \register[0][13] ,
         \register[0][12] , \register[0][11] , \register[0][10] ,
         \register[0][9] , \register[0][8] , \register[0][7] ,
         \register[0][6] , \register[0][5] , \register[0][4] ,
         \register[0][3] , \register[0][2] , \register[0][1] ,
         \register[0][0] , N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, n35, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287;
  wire   [1:0] fixedIndex;
  tri   [15:0] bus;

  TNBUFFHX1 \bus_tri[0]  ( .IN(N37), .ENB(rEn), .Q(bus[0]) );
  TNBUFFHX1 \bus_tri[1]  ( .IN(N36), .ENB(rEn), .Q(bus[1]) );
  TNBUFFHX1 \bus_tri[2]  ( .IN(N35), .ENB(rEn), .Q(bus[2]) );
  TNBUFFHX1 \bus_tri[3]  ( .IN(N34), .ENB(rEn), .Q(bus[3]) );
  TNBUFFHX1 \bus_tri[4]  ( .IN(N33), .ENB(rEn), .Q(bus[4]) );
  TNBUFFHX1 \bus_tri[5]  ( .IN(N32), .ENB(rEn), .Q(bus[5]) );
  TNBUFFHX1 \bus_tri[6]  ( .IN(N31), .ENB(rEn), .Q(bus[6]) );
  TNBUFFHX1 \bus_tri[7]  ( .IN(N30), .ENB(rEn), .Q(bus[7]) );
  TNBUFFHX1 \bus_tri[8]  ( .IN(N29), .ENB(rEn), .Q(bus[8]) );
  TNBUFFHX1 \bus_tri[9]  ( .IN(N28), .ENB(rEn), .Q(bus[9]) );
  TNBUFFHX1 \bus_tri[10]  ( .IN(N27), .ENB(rEn), .Q(bus[10]) );
  TNBUFFHX1 \bus_tri[11]  ( .IN(N26), .ENB(rEn), .Q(bus[11]) );
  TNBUFFHX1 \bus_tri[12]  ( .IN(N25), .ENB(rEn), .Q(bus[12]) );
  TNBUFFHX1 \bus_tri[13]  ( .IN(N24), .ENB(rEn), .Q(bus[13]) );
  TNBUFFHX1 \bus_tri[14]  ( .IN(N23), .ENB(rEn), .Q(bus[14]) );
  TNBUFFHX1 \bus_tri[15]  ( .IN(N22), .ENB(rEn), .Q(bus[15]) );
  DFFARX1 \register_reg[0][15]  ( .D(n124), .CLK(n278), .RSTB(n270), .Q(
        \register[0][15] ) );
  DFFARX1 \register_reg[0][14]  ( .D(n123), .CLK(n278), .RSTB(n270), .Q(
        \register[0][14] ) );
  DFFARX1 \register_reg[0][13]  ( .D(n122), .CLK(n278), .RSTB(n270), .Q(
        \register[0][13] ) );
  DFFARX1 \register_reg[0][12]  ( .D(n121), .CLK(n278), .RSTB(n270), .Q(
        \register[0][12] ) );
  DFFARX1 \register_reg[0][11]  ( .D(n120), .CLK(n278), .RSTB(n270), .Q(
        \register[0][11] ) );
  DFFARX1 \register_reg[0][10]  ( .D(n119), .CLK(n278), .RSTB(n270), .Q(
        \register[0][10] ) );
  DFFARX1 \register_reg[0][9]  ( .D(n118), .CLK(n278), .RSTB(n270), .Q(
        \register[0][9] ) );
  DFFARX1 \register_reg[0][8]  ( .D(n117), .CLK(n278), .RSTB(n269), .Q(
        \register[0][8] ) );
  DFFARX1 \register_reg[0][7]  ( .D(n116), .CLK(n277), .RSTB(n269), .Q(
        \register[0][7] ) );
  DFFARX1 \register_reg[0][6]  ( .D(n115), .CLK(n277), .RSTB(n269), .Q(
        \register[0][6] ) );
  DFFARX1 \register_reg[0][5]  ( .D(n114), .CLK(n277), .RSTB(n269), .Q(
        \register[0][5] ) );
  DFFARX1 \register_reg[0][4]  ( .D(n113), .CLK(n277), .RSTB(n269), .Q(
        \register[0][4] ) );
  DFFARX1 \register_reg[0][3]  ( .D(n112), .CLK(n277), .RSTB(n269), .Q(
        \register[0][3] ) );
  DFFARX1 \register_reg[0][2]  ( .D(n111), .CLK(n277), .RSTB(n269), .Q(
        \register[0][2] ) );
  DFFARX1 \register_reg[0][1]  ( .D(n110), .CLK(n277), .RSTB(n269), .Q(
        \register[0][1] ) );
  DFFARX1 \register_reg[0][0]  ( .D(n109), .CLK(n277), .RSTB(n269), .Q(
        \register[0][0] ) );
  DFFARX1 \register_reg[1][15]  ( .D(n140), .CLK(n280), .RSTB(n272), .Q(
        \register[1][15] ) );
  DFFARX1 \register_reg[1][14]  ( .D(n139), .CLK(n280), .RSTB(n272), .Q(
        \register[1][14] ) );
  DFFARX1 \register_reg[1][13]  ( .D(n138), .CLK(n280), .RSTB(n272), .Q(
        \register[1][13] ) );
  DFFARX1 \register_reg[1][12]  ( .D(n137), .CLK(n280), .RSTB(n272), .Q(
        \register[1][12] ) );
  DFFARX1 \register_reg[1][11]  ( .D(n136), .CLK(n280), .RSTB(n272), .Q(
        \register[1][11] ) );
  DFFARX1 \register_reg[1][10]  ( .D(n135), .CLK(n280), .RSTB(n271), .Q(
        \register[1][10] ) );
  DFFARX1 \register_reg[1][9]  ( .D(n134), .CLK(n280), .RSTB(n271), .Q(
        \register[1][9] ) );
  DFFARX1 \register_reg[1][8]  ( .D(n133), .CLK(n280), .RSTB(n271), .Q(
        \register[1][8] ) );
  DFFARX1 \register_reg[1][7]  ( .D(n132), .CLK(n279), .RSTB(n271), .Q(
        \register[1][7] ) );
  DFFARX1 \register_reg[1][6]  ( .D(n131), .CLK(n279), .RSTB(n271), .Q(
        \register[1][6] ) );
  DFFARX1 \register_reg[1][5]  ( .D(n130), .CLK(n279), .RSTB(n271), .Q(
        \register[1][5] ) );
  DFFARX1 \register_reg[1][4]  ( .D(n129), .CLK(n279), .RSTB(n271), .Q(
        \register[1][4] ) );
  DFFARX1 \register_reg[1][3]  ( .D(n128), .CLK(n279), .RSTB(n271), .Q(
        \register[1][3] ) );
  DFFARX1 \register_reg[1][2]  ( .D(n127), .CLK(n279), .RSTB(n271), .Q(
        \register[1][2] ) );
  DFFARX1 \register_reg[1][1]  ( .D(n126), .CLK(n279), .RSTB(n270), .Q(
        \register[1][1] ) );
  DFFARX1 \register_reg[1][0]  ( .D(n125), .CLK(n279), .RSTB(n270), .Q(
        \register[1][0] ) );
  DFFARX1 \register_reg[2][15]  ( .D(n156), .CLK(n282), .RSTB(n274), .Q(
        \register[2][15] ) );
  DFFARX1 \register_reg[2][14]  ( .D(n155), .CLK(n282), .RSTB(n274), .Q(
        \register[2][14] ) );
  DFFARX1 \register_reg[2][13]  ( .D(n154), .CLK(n282), .RSTB(n274), .Q(
        \register[2][13] ) );
  DFFARX1 \register_reg[2][12]  ( .D(n153), .CLK(n282), .RSTB(n273), .Q(
        \register[2][12] ) );
  DFFARX1 \register_reg[2][11]  ( .D(n152), .CLK(n282), .RSTB(n273), .Q(
        \register[2][11] ) );
  DFFARX1 \register_reg[2][10]  ( .D(n151), .CLK(n282), .RSTB(n273), .Q(
        \register[2][10] ) );
  DFFARX1 \register_reg[2][9]  ( .D(n150), .CLK(n282), .RSTB(n273), .Q(
        \register[2][9] ) );
  DFFARX1 \register_reg[2][8]  ( .D(n149), .CLK(n282), .RSTB(n273), .Q(
        \register[2][8] ) );
  DFFARX1 \register_reg[2][7]  ( .D(n148), .CLK(n281), .RSTB(n273), .Q(
        \register[2][7] ) );
  DFFARX1 \register_reg[2][6]  ( .D(n147), .CLK(n281), .RSTB(n273), .Q(
        \register[2][6] ) );
  DFFARX1 \register_reg[2][5]  ( .D(n146), .CLK(n281), .RSTB(n273), .Q(
        \register[2][5] ) );
  DFFARX1 \register_reg[2][4]  ( .D(n145), .CLK(n281), .RSTB(n273), .Q(
        \register[2][4] ) );
  DFFARX1 \register_reg[2][3]  ( .D(n144), .CLK(n281), .RSTB(n272), .Q(
        \register[2][3] ) );
  DFFARX1 \register_reg[2][2]  ( .D(n143), .CLK(n281), .RSTB(n272), .Q(
        \register[2][2] ) );
  DFFARX1 \register_reg[2][1]  ( .D(n142), .CLK(n281), .RSTB(n272), .Q(
        \register[2][1] ) );
  DFFARX1 \register_reg[2][0]  ( .D(n141), .CLK(n281), .RSTB(n272), .Q(
        \register[2][0] ) );
  DFFARX1 \register_reg[3][15]  ( .D(n172), .CLK(n284), .RSTB(n276), .Q(
        \register[3][15] ) );
  DFFARX1 \register_reg[3][14]  ( .D(n171), .CLK(n284), .RSTB(n275), .Q(
        \register[3][14] ) );
  DFFARX1 \register_reg[3][13]  ( .D(n170), .CLK(n284), .RSTB(n275), .Q(
        \register[3][13] ) );
  DFFARX1 \register_reg[3][12]  ( .D(n169), .CLK(n284), .RSTB(n275), .Q(
        \register[3][12] ) );
  DFFARX1 \register_reg[3][11]  ( .D(n168), .CLK(n284), .RSTB(n275), .Q(
        \register[3][11] ) );
  DFFARX1 \register_reg[3][10]  ( .D(n167), .CLK(n284), .RSTB(n275), .Q(
        \register[3][10] ) );
  DFFARX1 \register_reg[3][9]  ( .D(n166), .CLK(n284), .RSTB(n275), .Q(
        \register[3][9] ) );
  DFFARX1 \register_reg[3][8]  ( .D(n165), .CLK(n284), .RSTB(n275), .Q(
        \register[3][8] ) );
  DFFARX1 \register_reg[3][7]  ( .D(n164), .CLK(n283), .RSTB(n275), .Q(
        \register[3][7] ) );
  DFFARX1 \register_reg[3][6]  ( .D(n163), .CLK(n283), .RSTB(n275), .Q(
        \register[3][6] ) );
  DFFARX1 \register_reg[3][5]  ( .D(n162), .CLK(n283), .RSTB(n274), .Q(
        \register[3][5] ) );
  DFFARX1 \register_reg[3][4]  ( .D(n161), .CLK(n283), .RSTB(n274), .Q(
        \register[3][4] ) );
  DFFARX1 \register_reg[3][3]  ( .D(n160), .CLK(n283), .RSTB(n274), .Q(
        \register[3][3] ) );
  DFFARX1 \register_reg[3][2]  ( .D(n159), .CLK(n283), .RSTB(n274), .Q(
        \register[3][2] ) );
  DFFARX1 \register_reg[3][1]  ( .D(n158), .CLK(n283), .RSTB(n274), .Q(
        \register[3][1] ) );
  DFFARX1 \register_reg[3][0]  ( .D(n157), .CLK(n283), .RSTB(n274), .Q(
        \register[3][0] ) );
  DFFARX1 \fixedIndex_reg[1]  ( .D(index[1]), .CLK(rEn), .RSTB(n276), .Q(
        fixedIndex[1]) );
  DFFARX1 \fixedIndex_reg[0]  ( .D(index[0]), .CLK(rEn), .RSTB(n276), .Q(
        fixedIndex[0]) );
  NBUFFX2 U79 ( .IN(bus[0]), .Q(n175) );
  NBUFFX2 U80 ( .IN(bus[1]), .Q(n176) );
  NBUFFX2 U81 ( .IN(bus[2]), .Q(n177) );
  NBUFFX2 U82 ( .IN(bus[3]), .Q(n178) );
  NBUFFX2 U83 ( .IN(bus[4]), .Q(n179) );
  NBUFFX2 U84 ( .IN(bus[5]), .Q(n180) );
  NBUFFX2 U85 ( .IN(bus[6]), .Q(n181) );
  NBUFFX2 U86 ( .IN(bus[7]), .Q(n182) );
  NBUFFX2 U87 ( .IN(bus[8]), .Q(n183) );
  NBUFFX2 U88 ( .IN(bus[9]), .Q(n184) );
  NBUFFX2 U89 ( .IN(bus[10]), .Q(n185) );
  NBUFFX2 U90 ( .IN(bus[11]), .Q(n186) );
  NBUFFX2 U91 ( .IN(bus[12]), .Q(n187) );
  NBUFFX2 U92 ( .IN(bus[13]), .Q(n188) );
  NBUFFX2 U93 ( .IN(bus[14]), .Q(n189) );
  NBUFFX2 U94 ( .IN(bus[15]), .Q(n190) );
  INVX0 U95 ( .IN(n191), .QN(n262) );
  INVX0 U96 ( .IN(n191), .QN(n261) );
  AND3X1 U97 ( .IN1(n286), .IN2(n285), .IN3(n35), .Q(n191) );
  NBUFFX2 U98 ( .IN(n287), .Q(n269) );
  NBUFFX2 U99 ( .IN(n287), .Q(n270) );
  NBUFFX2 U100 ( .IN(n287), .Q(n271) );
  NBUFFX2 U101 ( .IN(n287), .Q(n272) );
  NBUFFX2 U102 ( .IN(n287), .Q(n273) );
  NBUFFX2 U103 ( .IN(n287), .Q(n274) );
  NBUFFX2 U104 ( .IN(n287), .Q(n275) );
  NBUFFX2 U105 ( .IN(n287), .Q(n276) );
  INVX0 U106 ( .IN(n192), .QN(n264) );
  INVX0 U107 ( .IN(n193), .QN(n266) );
  INVX0 U108 ( .IN(n194), .QN(n268) );
  INVX0 U109 ( .IN(n192), .QN(n263) );
  INVX0 U110 ( .IN(n193), .QN(n265) );
  INVX0 U111 ( .IN(n194), .QN(n267) );
  MUX41X1 U112 ( .IN1(\register[0][15] ), .IN3(\register[2][15] ), .IN2(
        \register[1][15] ), .IN4(\register[3][15] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N22) );
  MUX41X1 U113 ( .IN1(\register[0][14] ), .IN3(\register[2][14] ), .IN2(
        \register[1][14] ), .IN4(\register[3][14] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N23) );
  MUX41X1 U114 ( .IN1(\register[0][13] ), .IN3(\register[2][13] ), .IN2(
        \register[1][13] ), .IN4(\register[3][13] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N24) );
  MUX41X1 U115 ( .IN1(\register[0][12] ), .IN3(\register[2][12] ), .IN2(
        \register[1][12] ), .IN4(\register[3][12] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N25) );
  MUX41X1 U116 ( .IN1(\register[0][11] ), .IN3(\register[2][11] ), .IN2(
        \register[1][11] ), .IN4(\register[3][11] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N26) );
  MUX41X1 U117 ( .IN1(\register[0][10] ), .IN3(\register[2][10] ), .IN2(
        \register[1][10] ), .IN4(\register[3][10] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N27) );
  MUX41X1 U118 ( .IN1(\register[0][9] ), .IN3(\register[2][9] ), .IN2(
        \register[1][9] ), .IN4(\register[3][9] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N28) );
  MUX41X1 U119 ( .IN1(\register[0][8] ), .IN3(\register[2][8] ), .IN2(
        \register[1][8] ), .IN4(\register[3][8] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N29) );
  MUX41X1 U120 ( .IN1(\register[0][7] ), .IN3(\register[2][7] ), .IN2(
        \register[1][7] ), .IN4(\register[3][7] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N30) );
  MUX41X1 U121 ( .IN1(\register[0][6] ), .IN3(\register[2][6] ), .IN2(
        \register[1][6] ), .IN4(\register[3][6] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N31) );
  MUX41X1 U122 ( .IN1(\register[0][5] ), .IN3(\register[2][5] ), .IN2(
        \register[1][5] ), .IN4(\register[3][5] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N32) );
  MUX41X1 U123 ( .IN1(\register[0][4] ), .IN3(\register[2][4] ), .IN2(
        \register[1][4] ), .IN4(\register[3][4] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N33) );
  MUX41X1 U124 ( .IN1(\register[0][3] ), .IN3(\register[2][3] ), .IN2(
        \register[1][3] ), .IN4(\register[3][3] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N34) );
  MUX41X1 U125 ( .IN1(\register[0][2] ), .IN3(\register[2][2] ), .IN2(
        \register[1][2] ), .IN4(\register[3][2] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N35) );
  MUX41X1 U126 ( .IN1(\register[0][1] ), .IN3(\register[2][1] ), .IN2(
        \register[1][1] ), .IN4(\register[3][1] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N36) );
  MUX41X1 U127 ( .IN1(\register[0][0] ), .IN3(\register[2][0] ), .IN2(
        \register[1][0] ), .IN4(\register[3][0] ), .S0(fixedIndex[1]), .S1(
        fixedIndex[0]), .Q(N37) );
  NOR2X0 U128 ( .IN1(index[3]), .IN2(index[2]), .QN(n35) );
  AO22X1 U129 ( .IN1(n191), .IN2(n175), .IN3(\register[0][0] ), .IN4(n262), 
        .Q(n109) );
  AO22X1 U130 ( .IN1(n191), .IN2(n176), .IN3(\register[0][1] ), .IN4(n262), 
        .Q(n110) );
  AO22X1 U131 ( .IN1(n191), .IN2(n177), .IN3(\register[0][2] ), .IN4(n262), 
        .Q(n111) );
  AO22X1 U132 ( .IN1(n191), .IN2(n178), .IN3(\register[0][3] ), .IN4(n262), 
        .Q(n112) );
  AO22X1 U133 ( .IN1(n191), .IN2(n179), .IN3(\register[0][4] ), .IN4(n262), 
        .Q(n113) );
  AO22X1 U134 ( .IN1(n191), .IN2(n185), .IN3(\register[0][10] ), .IN4(n262), 
        .Q(n119) );
  AO22X1 U135 ( .IN1(n191), .IN2(n186), .IN3(\register[0][11] ), .IN4(n262), 
        .Q(n120) );
  AO22X1 U136 ( .IN1(n191), .IN2(n187), .IN3(\register[0][12] ), .IN4(n262), 
        .Q(n121) );
  AO22X1 U137 ( .IN1(n191), .IN2(n188), .IN3(\register[0][13] ), .IN4(n262), 
        .Q(n122) );
  AO22X1 U138 ( .IN1(n191), .IN2(n189), .IN3(\register[0][14] ), .IN4(n262), 
        .Q(n123) );
  AO22X1 U139 ( .IN1(n191), .IN2(n190), .IN3(\register[0][15] ), .IN4(n262), 
        .Q(n124) );
  AO22X1 U140 ( .IN1(n192), .IN2(n175), .IN3(\register[1][0] ), .IN4(n264), 
        .Q(n125) );
  AO22X1 U141 ( .IN1(n192), .IN2(n176), .IN3(\register[1][1] ), .IN4(n264), 
        .Q(n126) );
  AO22X1 U142 ( .IN1(n192), .IN2(n177), .IN3(\register[1][2] ), .IN4(n264), 
        .Q(n127) );
  AO22X1 U143 ( .IN1(n192), .IN2(n178), .IN3(\register[1][3] ), .IN4(n264), 
        .Q(n128) );
  AO22X1 U144 ( .IN1(n192), .IN2(n179), .IN3(\register[1][4] ), .IN4(n264), 
        .Q(n129) );
  AO22X1 U145 ( .IN1(n192), .IN2(n185), .IN3(\register[1][10] ), .IN4(n264), 
        .Q(n135) );
  AO22X1 U146 ( .IN1(n192), .IN2(n186), .IN3(\register[1][11] ), .IN4(n264), 
        .Q(n136) );
  AO22X1 U147 ( .IN1(n192), .IN2(n187), .IN3(\register[1][12] ), .IN4(n264), 
        .Q(n137) );
  AO22X1 U148 ( .IN1(n192), .IN2(n188), .IN3(\register[1][13] ), .IN4(n264), 
        .Q(n138) );
  AO22X1 U149 ( .IN1(n192), .IN2(n189), .IN3(\register[1][14] ), .IN4(n264), 
        .Q(n139) );
  AO22X1 U150 ( .IN1(n192), .IN2(n190), .IN3(\register[1][15] ), .IN4(n264), 
        .Q(n140) );
  AO22X1 U151 ( .IN1(n193), .IN2(n175), .IN3(\register[2][0] ), .IN4(n266), 
        .Q(n141) );
  AO22X1 U152 ( .IN1(n193), .IN2(n176), .IN3(\register[2][1] ), .IN4(n266), 
        .Q(n142) );
  AO22X1 U153 ( .IN1(n193), .IN2(n177), .IN3(\register[2][2] ), .IN4(n266), 
        .Q(n143) );
  AO22X1 U154 ( .IN1(n193), .IN2(n178), .IN3(\register[2][3] ), .IN4(n266), 
        .Q(n144) );
  AO22X1 U155 ( .IN1(n193), .IN2(n179), .IN3(\register[2][4] ), .IN4(n266), 
        .Q(n145) );
  AO22X1 U156 ( .IN1(n193), .IN2(n185), .IN3(\register[2][10] ), .IN4(n266), 
        .Q(n151) );
  AO22X1 U157 ( .IN1(n193), .IN2(n186), .IN3(\register[2][11] ), .IN4(n266), 
        .Q(n152) );
  AO22X1 U158 ( .IN1(n193), .IN2(n187), .IN3(\register[2][12] ), .IN4(n266), 
        .Q(n153) );
  AO22X1 U159 ( .IN1(n193), .IN2(n188), .IN3(\register[2][13] ), .IN4(n266), 
        .Q(n154) );
  AO22X1 U160 ( .IN1(n193), .IN2(n189), .IN3(\register[2][14] ), .IN4(n266), 
        .Q(n155) );
  AO22X1 U161 ( .IN1(n193), .IN2(n190), .IN3(\register[2][15] ), .IN4(n266), 
        .Q(n156) );
  AO22X1 U162 ( .IN1(n175), .IN2(n194), .IN3(\register[3][0] ), .IN4(n268), 
        .Q(n157) );
  AO22X1 U163 ( .IN1(n176), .IN2(n194), .IN3(\register[3][1] ), .IN4(n268), 
        .Q(n158) );
  AO22X1 U164 ( .IN1(n177), .IN2(n194), .IN3(\register[3][2] ), .IN4(n268), 
        .Q(n159) );
  AO22X1 U165 ( .IN1(n178), .IN2(n194), .IN3(\register[3][3] ), .IN4(n268), 
        .Q(n160) );
  AO22X1 U166 ( .IN1(n179), .IN2(n194), .IN3(\register[3][4] ), .IN4(n268), 
        .Q(n161) );
  AO22X1 U167 ( .IN1(n185), .IN2(n194), .IN3(\register[3][10] ), .IN4(n268), 
        .Q(n167) );
  AO22X1 U168 ( .IN1(n186), .IN2(n194), .IN3(\register[3][11] ), .IN4(n268), 
        .Q(n168) );
  AO22X1 U169 ( .IN1(n187), .IN2(n194), .IN3(\register[3][12] ), .IN4(n268), 
        .Q(n169) );
  AO22X1 U170 ( .IN1(n188), .IN2(n194), .IN3(\register[3][13] ), .IN4(n268), 
        .Q(n170) );
  AO22X1 U171 ( .IN1(n189), .IN2(n194), .IN3(\register[3][14] ), .IN4(n268), 
        .Q(n171) );
  AO22X1 U172 ( .IN1(n190), .IN2(n194), .IN3(\register[3][15] ), .IN4(n268), 
        .Q(n172) );
  AO22X1 U173 ( .IN1(n191), .IN2(n180), .IN3(\register[0][5] ), .IN4(n261), 
        .Q(n114) );
  AO22X1 U174 ( .IN1(n191), .IN2(n181), .IN3(\register[0][6] ), .IN4(n261), 
        .Q(n115) );
  AO22X1 U175 ( .IN1(n191), .IN2(n182), .IN3(\register[0][7] ), .IN4(n261), 
        .Q(n116) );
  AO22X1 U176 ( .IN1(n191), .IN2(n183), .IN3(\register[0][8] ), .IN4(n261), 
        .Q(n117) );
  AO22X1 U177 ( .IN1(n191), .IN2(n184), .IN3(\register[0][9] ), .IN4(n261), 
        .Q(n118) );
  AO22X1 U178 ( .IN1(n192), .IN2(n180), .IN3(\register[1][5] ), .IN4(n263), 
        .Q(n130) );
  AO22X1 U179 ( .IN1(n192), .IN2(n181), .IN3(\register[1][6] ), .IN4(n263), 
        .Q(n131) );
  AO22X1 U180 ( .IN1(n192), .IN2(n182), .IN3(\register[1][7] ), .IN4(n263), 
        .Q(n132) );
  AO22X1 U181 ( .IN1(n192), .IN2(n183), .IN3(\register[1][8] ), .IN4(n263), 
        .Q(n133) );
  AO22X1 U182 ( .IN1(n192), .IN2(n184), .IN3(\register[1][9] ), .IN4(n263), 
        .Q(n134) );
  AO22X1 U183 ( .IN1(n193), .IN2(n180), .IN3(\register[2][5] ), .IN4(n265), 
        .Q(n146) );
  AO22X1 U184 ( .IN1(n193), .IN2(n181), .IN3(\register[2][6] ), .IN4(n265), 
        .Q(n147) );
  AO22X1 U185 ( .IN1(n193), .IN2(n182), .IN3(\register[2][7] ), .IN4(n265), 
        .Q(n148) );
  AO22X1 U186 ( .IN1(n193), .IN2(n183), .IN3(\register[2][8] ), .IN4(n265), 
        .Q(n149) );
  AO22X1 U187 ( .IN1(n193), .IN2(n184), .IN3(\register[2][9] ), .IN4(n265), 
        .Q(n150) );
  AO22X1 U188 ( .IN1(n180), .IN2(n194), .IN3(\register[3][5] ), .IN4(n267), 
        .Q(n162) );
  AO22X1 U189 ( .IN1(n181), .IN2(n194), .IN3(\register[3][6] ), .IN4(n267), 
        .Q(n163) );
  AO22X1 U190 ( .IN1(n182), .IN2(n194), .IN3(\register[3][7] ), .IN4(n267), 
        .Q(n164) );
  AO22X1 U191 ( .IN1(n183), .IN2(n194), .IN3(\register[3][8] ), .IN4(n267), 
        .Q(n165) );
  AO22X1 U192 ( .IN1(n184), .IN2(n194), .IN3(\register[3][9] ), .IN4(n267), 
        .Q(n166) );
  AND3X1 U193 ( .IN1(n35), .IN2(n285), .IN3(index[0]), .Q(n192) );
  AND3X1 U194 ( .IN1(n35), .IN2(n286), .IN3(index[1]), .Q(n193) );
  AND3X1 U195 ( .IN1(index[0]), .IN2(n35), .IN3(index[1]), .Q(n194) );
  NBUFFX2 U196 ( .IN(wEn), .Q(n277) );
  NBUFFX2 U197 ( .IN(wEn), .Q(n278) );
  NBUFFX2 U198 ( .IN(wEn), .Q(n279) );
  NBUFFX2 U199 ( .IN(wEn), .Q(n280) );
  NBUFFX2 U200 ( .IN(wEn), .Q(n281) );
  NBUFFX2 U201 ( .IN(wEn), .Q(n282) );
  NBUFFX2 U202 ( .IN(wEn), .Q(n283) );
  NBUFFX2 U203 ( .IN(wEn), .Q(n284) );
  INVX0 U204 ( .IN(reset), .QN(n287) );
  INVX0 U205 ( .IN(index[1]), .QN(n285) );
  INVX0 U206 ( .IN(index[0]), .QN(n286) );
endmodule

